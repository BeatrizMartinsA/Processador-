module add(entrada1, entrada2, saida);
input [31:0] entrada1, entrada2;
output [31:0] saida;

assign saida = entrada1 + entrada2;

endmodule
